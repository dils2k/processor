module lab00_test(
  input clk,
  output clk1
);

assign clk1 = clk;

endmodule
